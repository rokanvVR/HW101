`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.10.2025 21:18:27
// Design Name: 
// Module Name: wires4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module wires4(
    input a,b,c,
    input w,x,y,z
    );
    assign w =a;
    assign x = b;
    assign y = b;
    assign z = c;
endmodule
